module bluemux(I,inA,inB,outA,outB)
    


endmodule 