//Spencer Dugas
//Andrew Doucet

//Move to move contents of register A to register B

module MOV (RA, RB);
    input [15:0] RA;
    output [15:0] RB;

    assign RB = RA;
    
endmodule
    
